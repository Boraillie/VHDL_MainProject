library verilog;
use verilog.vl_types.all;
entity fulladder_nbitsand_N4_1 is
    port(
        sin_i           : in     vl_logic_vector(3 downto 0);
        op1_i           : in     vl_logic_vector(3 downto 0);
        op2j_i          : in     vl_logic;
        cin_i           : in     vl_logic;
        s_o             : out    vl_logic_vector(3 downto 0);
        cout_o          : out    vl_logic
    );
end fulladder_nbitsand_N4_1;
